module gate_xor(input x, y,output z);
	xor(z, x, y);
endmodule

module gate_and(input x, y,output z);
	and(z, x, y);
endmodule

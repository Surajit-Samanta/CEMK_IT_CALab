module gate_or(input x, y,output z);
	or(z, x, y);
endmodule

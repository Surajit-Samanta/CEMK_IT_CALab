module gate_nand(input x, y,output z);
	nand(z, x, y);
endmodule

module gate_nor(input x, y,output z);
	nor(z, x, y);
endmodule

module gate_xnor(input x, y,output z);
	xnor(z, x, y);
endmodule

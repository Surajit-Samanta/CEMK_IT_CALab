module hello;
 initial
	begin
		$display("Name:- Surajit Samanta\nRoll no:- IT\23\L69\nDept:- Information Technology\nSem:- 4th");
		$finish;
	end
endmodule	
